module table

pub fn say() {
	println('helle')
}